module half_adder( 
    input a, b,
    output cout, sum );
	
    assign {cout, sum} = a + b;
endmodule